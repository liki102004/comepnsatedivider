module LED2(a,b);

input [7:0] a; //피제수 
output reg b;//signal

always@(a or b)
begin
if(a==35||a==39||
	a==43||a==47||
	a==51||a==55||
	a==59||a==63||//4간격 ->2bit

	a==69||a==70||a==71||
	a==77||a==78||a==79||
	a==85||a==86||a==87||
	a==93||a==94||a==95||
	a==101||a==102||a==103||
	a==109||a==110||a==111||
	a==117||a==118||a==119||
	a==125||a==126||a==127||//8간격->3bit11
	
	a==137||a==138||a==139||a==140||a==141||a==142||a==143||
	a==153||a==154||a==155||a==156||a==157||a==158||a==159||
	a==169||a==170||a==171||a==172||a==173||a==174||a==175||
	a==185||a==186||a==187||a==188||a==189||a==190||a==191||
	a==201||a==202||a==203||a==204||a==205||a==206||a==207||
	a==217||a==218||a==219||a==220||a==221||a==222||a==223||
	//
	a==233||a==234||a==235||a==236||a==237||a==238||a==239||
	a==249||a==250||a==251||a==252||a==253||a==254||a==255)//16간격 
	b=1;
else
	b=0;
end
endmodule


